`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:35:30 06/03/2012 
// Design Name: 
// Module Name:    generarCircunferencia 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module generarCircunferencia(circunferencia);

output reg [15:0] circunferencia;
initial begin 

circunferencia = 2326;

end

endmodule
