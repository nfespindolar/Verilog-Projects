`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   13:40:14 05/15/2012
// Design Name:   vga_sync
// Module Name:   C:/Users/Fernando/Desktop/SimulacionesX/PrimerVGA/TestVGAsync.v
// Project Name:  PrimerVGA
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: vga_sync
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module TestVGAsync;

	// Outputs
	wire ;

	// Instantiate the Unit Under Test (UUT)
	vga_sync uut (
		.()
	);

	initial begin
		// Initialize Inputs

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
      
endmodule

